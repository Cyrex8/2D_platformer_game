    ����          Assembly-CSharp   Saver+Position   xyz      �@LR�� ��=